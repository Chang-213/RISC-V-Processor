module mp3_tb;
`timescale 1ns/10ps

/********************* Do not touch for proper compilation *******************/
// Instantiate Interfaces
tb_itf itf();
rvfi_itf rvfi(itf.clk, itf.rst);

// Instantiate Testbench
source_tb tb(
    .magic_mem_itf(itf),
    .mem_itf(itf),
    .sm_itf(itf),
    .tb_itf(itf),
    .rvfi(rvfi)
);
/****************************** End do not touch *****************************/
logic clk;
assign clk = itf.clk;
/************************ Signals necessary for monitor **********************/
// This section not required until CP3

assign rvfi.commit = 0; // Set high when a valid instruction is modifying regfile or PC
// Set high when you detect an infinite loop
assign rvfi.halt = dut.datapath.load_pc & ((dut.datapath.pc_out + 20) == dut.datapath.pc_d_out);
initial rvfi.order = 0;
always @(posedge itf.clk iff rvfi.commit) rvfi.order <= rvfi.order + 1; // Modify for OoO
/**************************** End RVFIMON signals ****************************/

/********************* Assign Shadow Memory Signals Here *********************/
// This section not required until CP2
/*********************** End Shadow Memory Assignments ***********************/

// Set this to the proper value
assign itf.registers = dut.datapath.regfile.data;

/*********************** Instantiate your design here ************************/
mp3 dut(
	.clk 			 (itf.clk),
	.rst 			 (itf.rst),
	.inst_resp		 (itf.inst_resp),
	.inst_rdata		 (itf.inst_rdata),
	.data_resp		 (itf.data_resp),
	.data_rdata		 (itf.data_rdata),
	.inst_read		 (itf.inst_read),
	.inst_addr		 (itf.inst_addr),
	.data_read		 (itf.data_read),
	.data_write		 (itf.data_write),
	.data_mbe		 (itf.data_mbe),
	.data_addr		 (itf.data_addr),
	.data_wdata		 (itf.data_wdata)
);
/***************************** End Instantiation *****************************/

endmodule
